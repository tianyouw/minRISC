// sys_pll.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module sys_pll (
		input  wire  ref_clk_clk,        //      ref_clk.clk
		input  wire  ref_reset_reset,    //    ref_reset.reset
		output wire  reset_source_reset, // reset_source.reset
		output wire  sdram_clk_clk,      //    sdram_clk.clk
		output wire  sys_clk_clk         //      sys_clk.clk
	);

	sys_pll_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),      //    sdram_clk.clk
		.reset_source_reset (reset_source_reset)  // reset_source.reset
	);

endmodule
